module AddSum(InA,InB,Result);

input [31:0] InA;
input [31:0] InB;

output [31:0] Result;

assign Result = InA + InB;




endmodule
