module ROM(out,address);

output reg [31:0] out;

input [31:0] address;


always @(address) begin
//00000203
	case (address)
	32'h00: out <= 32'h00400093; //addi 1
	32'h04: out <= 32'h00800113; // addi2
	32'h08: out <= 32'h002081B3;//Add
	32'h0c: out <= 32'h00100023; // store 1
	32'h10: out <= 32'h00200223; // Store 2
	32'h14: out <= 32'h00000203; // Load 1
	32'h18: out <= 32'h40210463; // beq
	
  // 8'h00: out <= 32'h00450693;//0000000 00100 01010 000 01101 0010011
  // 8'h04: out <= 32'h00100713;//0000000 00001 00000 000 01110 0010011
  // 8'h08: out <= 32'h00b76463;//0000000 01011 01110 110 01000 1100011
  // 8'h0c: out <= 32'h00008067;//0000000 00000 00001 000 00000 1100111
  // 8'h10: out <= 32'h0006a803;//0000000 00000 01101 010 10000 0000011
  // 8'h14: out <= 32'h00068613;//0000000 00000 01101 000 01100 0010011
  // 8'h18: out <= 32'h00070793;//0000000 00000 01110 000 01111 0010011
  // 8'h1c: out <= 32'hffc62883;//1111111 11100 01100 010 10001 0000011
  // 8'h20: out <= 32'h01185a63;//0000000 10001 10000 101 10100 1100011
   //8'h24: out <= 32'h01162023;//0000000 10001 01100 010 00000 0100011
   //8'h28: out <= 32'hfff78793;//1111111 11111 01111 000 01111 0010011
   //8'h2c: out <= 32'hffc60613;//1111111 11100 01100 000 01100 0010011
  // 8'h30: out <= 32'hfe0796e3;//1111111 00000 01111 001 01101 1100011
  // 8'h34: out <= 32'h00279793;//0000000 00010 01111 001 01111 0010011
   //8'h38: out <= 32'h00f507b3;//0000000 01111 01010 000 01111 0110011
   //8'h3c: out <= 32'h0107a023;//0000000 10000 01111 010 00000 0100011
   //8'h40: out <= 32'h00170713;//0000000 00001 01110 000 01110 0010011
   //8'h44: out <= 32'h00468693;//0000000 00100 01101 000 01101 0010011
   //8'h48: out <= 32'hfc1ff06f;//1111110 00001 11111 111 00000 1101111
	default: out <= 32'hxxxxxxxx;// nothing


endcase

end

endmodule